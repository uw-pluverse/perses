module test;

  // Thread gets started at the beginning of the simulation
  initial begin

    // Call to system task to print output in simulator console
    $display("Hello world!");
  end

endmodule