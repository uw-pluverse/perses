




module t;
   reg foobar;

   task boobar; endtask

   initial begin
      if (foobat) $stop;
      boobat;
   end
endmodule
