module test;
  initial
     display("Hello world!");
endmodule
