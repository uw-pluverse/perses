module t ;
reg foobar ;
task boobar ; endtask
initial begin
if ( boobar ) $ stop ;
boobat ;
end
endmodule
