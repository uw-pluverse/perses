

`define wxyz
